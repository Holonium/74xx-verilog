module mod_7405 (
	input A1, output Y1,
	input A2, output Y2,
	input A3, output Y3,
	input A4, output Y4,
	input A5, output Y5,
	input A6, output Y6
);
	assign Y1 = !A1;
	assign Y2 = !A2;
	assign Y3 = !A3;
	assign Y4 = !A4;
	assign Y5 = !A5;
	assign Y6 = !A6;
endmodule
