module mod_7430 (
	input A1, input B1, input C1, input D1, input E1, input F1, input G1, input H1, output Y1
);
	assign Y1 = !(A1 & B1 & C1 & D1 & E1 & F1 & G1 & H1);
endmodule
